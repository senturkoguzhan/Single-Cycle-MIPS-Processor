`define DELAY 20
module ALU_32BIT_testbench(); 
    wire [31:0]resAlu32;
    wire c_out;
	 wire V;
	 wire Z;
    reg [31:0]A;
    reg [31:0]B;
    reg [2:0]OP;

ALU_32BIT alu32tb(resAlu32,c_out,V,Z,A,B,OP);

initial begin
A = 32'b10101010101010101010101010101010; 
B = 32'b01010101010101010101010101010101;
OP = 3'b000;
#`DELAY;
A = 32'b10101010101010101010101010101010; 
B = 32'b01010101010101010101010101010101;
OP = 3'b001;
#`DELAY;
A = 32'b00000000000000000000000000001100; 
B = 32'b00000000000000000000000000001010;
OP = 3'b010;
#`DELAY;
A = 32'b00000000000000000000000000001100; 
B = 32'b00000000000000000000000000001010;
OP = 3'b110;
#`DELAY;
A = 32'b00000000000000000000000000001100; 
B = 32'b00000000000000000000000000001100;
OP = 3'b110;
#`DELAY;
A = 32'b11111111111111111111111111111111; 
B = 32'b11111111111111111111111111111111;
OP = 3'b010;
#`DELAY;
B = 32'b11111111111111111111111111111111; 
A = 32'b00000000000000000000000000000000;
OP = 3'b111;
end
 
 
initial
begin
$monitor("time = %2d, A =%32b, B =%32b, OP =%3b, R =%32b c_out =%1b Z=%1b", $time, A, B, OP ,resAlu32,c_out, Z);
end
 
endmodule