`define DELAY 20
module MUX_8X1_32_testbench(); 

	wire [31:0] out;
	reg [31:0] a1;
	reg [31:0] a2;
	reg [31:0] a3;
	reg [31:0] a4;
	reg [31:0] a5;
	reg [31:0] a6;
	reg [31:0] a7;
	reg [31:0] a8;
	reg [2:0] s;
	
MUX_8X1_32 mux8x132tb(out, a1,a2,a3,a4,a5,a6,a7,a8,s);

initial begin
a1 = 32'h00000000;
a2 = 32'h00000001;
a3 = 32'h00000002;
a4 = 32'h00000003;
a5 = 32'h00000004;
a6 = 32'h00000005;
a7 = 32'h00000006;
a8 = 32'h00000007;
s = 3'b000;
#`DELAY;
a1 = 32'h00000000;
a2 = 32'h00000001;
a3 = 32'h00000002;
a4 = 32'h00000003;
a5 = 32'h00000004;
a6 = 32'h00000005;
a7 = 32'h00000006;
a8 = 32'h00000007;
s = 3'b001;
#`DELAY;
a1 = 32'h00000000;
a2 = 32'h00000001;
a3 = 32'h00000002;
a4 = 32'h00000003;
a5 = 32'h00000004;
a6 = 32'h00000005;
a7 = 32'h00000006;
a8 = 32'h00000007;
s = 3'b10;
#`DELAY;
a1 = 32'h00000000;
a2 = 32'h00000001;
a3 = 32'h00000002;
a4 = 32'h00000003;
a5 = 32'h00000004;
a6 = 32'h00000005;
a7 = 32'h00000006;
a8 = 32'h00000007;
s = 3'b011;
#`DELAY;
a1 = 32'h00000000;
a2 = 32'h00000001;
a3 = 32'h00000002;
a4 = 32'h00000003;
a5 = 32'h00000004;
a6 = 32'h00000005;
a7 = 32'h00000006;
a8 = 32'h00000007;
s = 3'b100;
#`DELAY;
a1 = 32'h00000000;
a2 = 32'h00000001;
a3 = 32'h00000002;
a4 = 32'h00000003;
a5 = 32'h00000004;
a6 = 32'h00000005;
a7 = 32'h00000006;
a8 = 32'h00000007;
s = 3'b101;
#`DELAY;
a1 = 32'h00000000;
a2 = 32'h00000001;
a3 = 32'h00000002;
a4 = 32'h00000003;
a5 = 32'h00000004;
a6 = 32'h00000005;
a7 = 32'h00000006;
a8 = 32'h00000007;
s = 3'b110;
#`DELAY;
a1 = 32'h00000000;
a2 = 32'h00000001;
a3 = 32'h00000002;
a4 = 32'h00000003;
a5 = 32'h00000004;
a6 = 32'h00000005;
a7 = 32'h00000006;
a8 = 32'h00000007;
s = 3'b111;
#`DELAY;

end
 
initial
begin
$monitor("a1 =%32b, a2=%32b, a3=%32b ,a4=%32b ,a5 =%32b, a6=%32b, a7=%32b ,a8=%32b, s=%3b ,out=%32b ", a1,a2,a3,a4,a5,a6,a7,a8,s, out);
end
 
endmodule